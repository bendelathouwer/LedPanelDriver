module test1 (
    output R0in ,
    //output B0in ,
    output R1in ,
    //output B1in ,
    //output A0in ,
    //output A2in ,
    output SCLKin ,
    output BLANKin ,
    //output G0in ,
    //output G1in ,
    //output A4in ,
    //output A1in ,
    //output A3in,
    output LATCHin
);

reg [63:0] data ;

